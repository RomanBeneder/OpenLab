-- MC8051 IP Core Demo Design, Configuration for Top-level Design
-- Date: 2013-02-25
-- http://embsys.technikum-wien.at

configuration fpga_top_rtl_cfg of fpga_top is
    for rtl
    end for;
end fpga_top_rtl_cfg;
