-- MC8051 IP Core Demo Design, Configuration for Top-level Testbench 
-- Date: 2013-02-25
-- http://embsys.technikum-wien.at

configuration testbench_sim_cfg of testbench is
  for sim
  end for;
end testbench_sim_cfg;
