-- MC8051 IP Core Demo Design, Entity for Top-level Testbench 
-- Date: 2013-02-25
-- http://embsys.technikum-wien.at

library ieee;
use ieee.std_logic_1164.all;

use std.textio.all;

entity testbench is
end;
